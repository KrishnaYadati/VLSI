`timescale 1ns / 1ps
module HA(a,b,c,diff,borrow);
input a,b,c; output diff,borrow;
assign diff=a^b^c;
assign borrow=((~a)&b)|(b&c)|(c&(~a));
endmodule
